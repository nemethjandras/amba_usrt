//shift reg module

module 
